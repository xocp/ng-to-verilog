module ZERO16(
	output [15:0] OUT
);

assign OUT = 0;

endmodule
