module mraddressbus(
	output [15:0] OUT0,
	input [15:0] SRC,
	input [15:0] PC,
	input [15:0] AH_ACC,
	input [15:0] PG0_IDX0,
	input [15:0] PG1_IDX1
);

wire SPLIT16_0_D15;
wire SPLIT16_0_D14;
wire SPLIT16_0_D13;
wire SPLIT16_0_D12;
wire SPLIT16_0_D11;
wire SPLIT16_0_D10;
wire SPLIT16_0_D9;
wire SPLIT16_0_D8;
wire SPLIT16_0_D7;
wire SPLIT16_0_D6;
wire SPLIT16_0_D5;
wire SPLIT16_0_D4;
wire SPLIT16_0_D3;
wire SPLIT16_0_D2;
wire SPLIT16_0_D1;
wire SPLIT16_0_D0;
wire [15:0] SELECT16_1_OUT;
wire [15:0] SELECT16_2_OUT;
wire [15:0] SELECT16_3_OUT;
wire [15:0] ZERO16_4_OUT;
wire [15:0] SELECT16_5_OUT;

SPLIT16 SPLIT16_0(
	.D15 (SPLIT16_0_D15),
	.D14 (SPLIT16_0_D14),
	.D13 (SPLIT16_0_D13),
	.D12 (SPLIT16_0_D12),
	.D11 (SPLIT16_0_D11),
	.D10 (SPLIT16_0_D10),
	.D9 (SPLIT16_0_D9),
	.D8 (SPLIT16_0_D8),
	.D7 (SPLIT16_0_D7),
	.D6 (SPLIT16_0_D6),
	.D5 (SPLIT16_0_D5),
	.D4 (SPLIT16_0_D4),
	.D3 (SPLIT16_0_D3),
	.D2 (SPLIT16_0_D2),
	.D1 (SPLIT16_0_D1),
	.D0 (SPLIT16_0_D0),
	.IN (SRC)
);
	
SELECT16 SELECT16_1(
	.OUT (SELECT16_1_OUT),
	.S (SPLIT16_0_D4),
	.D1 (SELECT16_3_OUT),
	.D0 (SELECT16_2_OUT)
);
	
SELECT16 SELECT16_2(
	.OUT (SELECT16_2_OUT),
	.S (SPLIT16_0_D3),
	.D1 (AH_ACC),
	.D0 (PC)
);
	
SELECT16 SELECT16_3(
	.OUT (SELECT16_3_OUT),
	.S (SPLIT16_0_D3),
	.D1 (PG1_IDX1),
	.D0 (PG0_IDX0)
);
	
ZERO16 ZERO16_4(
	.OUT (ZERO16_4_OUT)
);
	
SELECT16 SELECT16_5(
	.OUT (SELECT16_5_OUT),
	.S (SPLIT16_0_D7),
	.D1 (SELECT16_1_OUT),
	.D0 (ZERO16_4_OUT)
);
	
assign OUT0 = SELECT16_5_OUT;

endmodule
