module ZERO(
	output OUT
);

assign OUT = 0;

endmodule
