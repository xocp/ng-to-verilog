module INC16(
	output [15:0] OUT,
	input [15:0] IN
);

assign OUT = IN + 1;

endmodule
