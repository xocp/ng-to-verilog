module NAND(
	output OUT,
	input A,
	input B
);

nand(OUT,A,B);

endmodule
