module mrspregister(
	output [15:0] HI,
	output [15:0] LO,
	output [15:0] HI_LO,
	input [15:0] D_IN,
	input A0,
	input STO,
	input STO_A,
	input [15:0] A_IN,
	input CLK
);

wire [15:0] DFF16_0_OUT;
wire [15:0] BUNDLE16_1_OUT;
wire [15:0] BUNDLE16_2_OUT;
wire SPLIT16_3_D15;
wire SPLIT16_3_D14;
wire SPLIT16_3_D13;
wire SPLIT16_3_D12;
wire SPLIT16_3_D11;
wire SPLIT16_3_D10;
wire SPLIT16_3_D9;
wire SPLIT16_3_D8;
wire SPLIT16_3_D7;
wire SPLIT16_3_D6;
wire SPLIT16_3_D5;
wire SPLIT16_3_D4;
wire SPLIT16_3_D3;
wire SPLIT16_3_D2;
wire SPLIT16_3_D1;
wire SPLIT16_3_D0;
wire OR_4_OUT;
wire SPLIT16_5_D15;
wire SPLIT16_5_D14;
wire SPLIT16_5_D13;
wire SPLIT16_5_D12;
wire SPLIT16_5_D11;
wire SPLIT16_5_D10;
wire SPLIT16_5_D9;
wire SPLIT16_5_D8;
wire SPLIT16_5_D7;
wire SPLIT16_5_D6;
wire SPLIT16_5_D5;
wire SPLIT16_5_D4;
wire SPLIT16_5_D3;
wire SPLIT16_5_D2;
wire SPLIT16_5_D1;
wire SPLIT16_5_D0;
wire SPLIT22_6_D21;
wire SPLIT22_6_D20;
wire SPLIT22_6_D19;
wire SPLIT22_6_D18;
wire SPLIT22_6_D17;
wire SPLIT22_6_D16;
wire SPLIT22_6_D15;
wire SPLIT22_6_D14;
wire SPLIT22_6_D13;
wire SPLIT22_6_D12;
wire SPLIT22_6_D11;
wire SPLIT22_6_D10;
wire SPLIT22_6_D9;
wire SPLIT22_6_D8;
wire SPLIT22_6_D7;
wire SPLIT22_6_D6;
wire SPLIT22_6_D5;
wire SPLIT22_6_D4;
wire SPLIT22_6_D3;
wire SPLIT22_6_D2;
wire SPLIT22_6_D1;
wire SPLIT22_6_D0;
wire [15:0] BUNDLE16_7_OUT;
wire [15:0] BUNDLE16_8_OUT;
wire [15:0] SELECT16_9_OUT;
wire [15:0] SELECT16_10_OUT;
wire ZERO_11_OUT;
wire ZERO_12_OUT;

DFF16 DFF16_0(
	.OUT (DFF16_0_OUT),
	.ST (OR_4_OUT),
	.X (SELECT16_10_OUT),
	.CLK (CLK)
);
	
BUNDLE16 BUNDLE16_1(
	.OUT (BUNDLE16_1_OUT),
	.D15 (ZERO_11_OUT),
	.D14 (ZERO_11_OUT),
	.D13 (ZERO_11_OUT),
	.D12 (ZERO_11_OUT),
	.D11 (ZERO_11_OUT),
	.D10 (ZERO_11_OUT),
	.D9 (ZERO_11_OUT),
	.D8 (ZERO_11_OUT),
	.D7 (SPLIT16_3_D15),
	.D6 (SPLIT16_3_D14),
	.D5 (SPLIT16_3_D13),
	.D4 (SPLIT16_3_D12),
	.D3 (SPLIT16_3_D11),
	.D2 (SPLIT16_3_D10),
	.D1 (SPLIT16_3_D9),
	.D0 (SPLIT16_3_D8)
);
	
BUNDLE16 BUNDLE16_2(
	.OUT (BUNDLE16_2_OUT),
	.D15 (ZERO_12_OUT),
	.D14 (ZERO_12_OUT),
	.D13 (ZERO_12_OUT),
	.D12 (ZERO_12_OUT),
	.D11 (ZERO_12_OUT),
	.D10 (ZERO_12_OUT),
	.D9 (ZERO_12_OUT),
	.D8 (ZERO_12_OUT),
	.D7 (SPLIT16_3_D7),
	.D6 (SPLIT16_3_D6),
	.D5 (SPLIT16_3_D5),
	.D4 (SPLIT16_3_D4),
	.D3 (SPLIT16_3_D3),
	.D2 (SPLIT16_3_D2),
	.D1 (SPLIT16_3_D1),
	.D0 (SPLIT16_3_D0)
);
	
SPLIT16 SPLIT16_3(
	.D15 (SPLIT16_3_D15),
	.D14 (SPLIT16_3_D14),
	.D13 (SPLIT16_3_D13),
	.D12 (SPLIT16_3_D12),
	.D11 (SPLIT16_3_D11),
	.D10 (SPLIT16_3_D10),
	.D9 (SPLIT16_3_D9),
	.D8 (SPLIT16_3_D8),
	.D7 (SPLIT16_3_D7),
	.D6 (SPLIT16_3_D6),
	.D5 (SPLIT16_3_D5),
	.D4 (SPLIT16_3_D4),
	.D3 (SPLIT16_3_D3),
	.D2 (SPLIT16_3_D2),
	.D1 (SPLIT16_3_D1),
	.D0 (SPLIT16_3_D0),
	.IN (DFF16_0_OUT)
);
	
OR OR_4(
	.OUT (OR_4_OUT),
	.A (STO),
	.B (STO_A)
);
	
SPLIT16 SPLIT16_5(
	.D15 (SPLIT16_5_D15),
	.D14 (SPLIT16_5_D14),
	.D13 (SPLIT16_5_D13),
	.D12 (SPLIT16_5_D12),
	.D11 (SPLIT16_5_D11),
	.D10 (SPLIT16_5_D10),
	.D9 (SPLIT16_5_D9),
	.D8 (SPLIT16_5_D8),
	.D7 (SPLIT16_5_D7),
	.D6 (SPLIT16_5_D6),
	.D5 (SPLIT16_5_D5),
	.D4 (SPLIT16_5_D4),
	.D3 (SPLIT16_5_D3),
	.D2 (SPLIT16_5_D2),
	.D1 (SPLIT16_5_D1),
	.D0 (SPLIT16_5_D0),
	.IN (D_IN)
);
	
SPLIT22 SPLIT22_6(
	.D21 (SPLIT22_6_D21),
	.D20 (SPLIT22_6_D20),
	.D19 (SPLIT22_6_D19),
	.D18 (SPLIT22_6_D18),
	.D17 (SPLIT22_6_D17),
	.D16 (SPLIT22_6_D16),
	.D15 (SPLIT22_6_D15),
	.D14 (SPLIT22_6_D14),
	.D13 (SPLIT22_6_D13),
	.D12 (SPLIT22_6_D12),
	.D11 (SPLIT22_6_D11),
	.D10 (SPLIT22_6_D10),
	.D9 (SPLIT22_6_D9),
	.D8 (SPLIT22_6_D8),
	.D7 (SPLIT22_6_D7),
	.D6 (SPLIT22_6_D6),
	.D5 (SPLIT22_6_D5),
	.D4 (SPLIT22_6_D4),
	.D3 (SPLIT22_6_D3),
	.D2 (SPLIT22_6_D2),
	.D1 (SPLIT22_6_D1),
	.D0 (SPLIT22_6_D0),
	.IN (DFF16_0_OUT)
);
	
BUNDLE16 BUNDLE16_7(
	.OUT (BUNDLE16_7_OUT),
	.D15 (SPLIT16_5_D7),
	.D14 (SPLIT16_5_D6),
	.D13 (SPLIT16_5_D5),
	.D12 (SPLIT16_5_D4),
	.D11 (SPLIT16_5_D3),
	.D10 (SPLIT16_5_D2),
	.D9 (SPLIT16_5_D1),
	.D8 (SPLIT16_5_D0),
	.D7 (SPLIT22_6_D7),
	.D6 (SPLIT22_6_D6),
	.D5 (SPLIT22_6_D5),
	.D4 (SPLIT22_6_D4),
	.D3 (SPLIT22_6_D3),
	.D2 (SPLIT22_6_D2),
	.D1 (SPLIT22_6_D1),
	.D0 (SPLIT22_6_D0)
);
	
BUNDLE16 BUNDLE16_8(
	.OUT (BUNDLE16_8_OUT),
	.D15 (SPLIT22_6_D15),
	.D14 (SPLIT22_6_D14),
	.D13 (SPLIT22_6_D13),
	.D12 (SPLIT22_6_D12),
	.D11 (SPLIT22_6_D11),
	.D10 (SPLIT22_6_D10),
	.D9 (SPLIT22_6_D9),
	.D8 (SPLIT22_6_D8),
	.D7 (SPLIT16_5_D7),
	.D6 (SPLIT16_5_D6),
	.D5 (SPLIT16_5_D5),
	.D4 (SPLIT16_5_D4),
	.D3 (SPLIT16_5_D3),
	.D2 (SPLIT16_5_D2),
	.D1 (SPLIT16_5_D1),
	.D0 (SPLIT16_5_D0)
);
	
SELECT16 SELECT16_9(
	.OUT (SELECT16_9_OUT),
	.S (A0),
	.D1 (BUNDLE16_7_OUT),
	.D0 (BUNDLE16_8_OUT)
);
	
SELECT16 SELECT16_10(
	.OUT (SELECT16_10_OUT),
	.S (STO_A),
	.D1 (A_IN),
	.D0 (SELECT16_9_OUT)
);
	
ZERO ZERO_11(
	.OUT (ZERO_11_OUT)
);
	
ZERO ZERO_12(
	.OUT (ZERO_12_OUT)
);
	
assign HI = BUNDLE16_1_OUT;
assign LO = BUNDLE16_2_OUT;
assign HI_LO = DFF16_0_OUT;

endmodule
