module XOR16(
	output [15:0] OUT,
	input [15:0] A,
	input [15:0] B
);

assign OUT = A ^ B;

endmodule
